library verilog;
use verilog.vl_types.all;
entity test_padder1 is
end test_padder1;
