library verilog;
use verilog.vl_types.all;
entity tb_iota is
end tb_iota;
