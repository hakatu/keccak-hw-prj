library verilog;
use verilog.vl_types.all;
entity test_padder is
end test_padder;
