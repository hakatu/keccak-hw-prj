library verilog;
use verilog.vl_types.all;
entity tb_keccak_round is
end tb_keccak_round;
