library verilog;
use verilog.vl_types.all;
entity test_keccak is
end test_keccak;
