library verilog;
use verilog.vl_types.all;
entity keccak_f_1600_tb is
end keccak_f_1600_tb;
