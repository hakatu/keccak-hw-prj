library verilog;
use verilog.vl_types.all;
entity test_rconst2in1 is
end test_rconst2in1;
