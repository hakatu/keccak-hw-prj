library verilog;
use verilog.vl_types.all;
entity test_f_permutation is
end test_f_permutation;
