/* Keccak Core
	Module: string to array
	Date: 31/12/2021
	Author: Tran Cong Tien
	ID: 1810580
*/
import keccak_pkg::plane;
import keccak_pkg::state;
import keccak_pkg::N;

module string_to_array(s,a);
	input	[1599:0] s;
	output	state	 a;

always_comb
begin
	/*
	a[0][0] = {s[63:56], s[55:48], s[47:40], s[39:32], s[31:24], s[23:16], s[15:8], s[7:0]};
	a[0][1] = {s[127:120], s[119:112], s[111:104], s[103:96], s[95:88], s[87:80], s[79:72], s[71:64]};
	a[0][2] = {s[191:184], s[183:176], s[175:168], s[167:160], s[159:152], s[151:144], s[143:136], s[135:128]};
	a[0][3] = {s[255:248], s[247:240], s[239:232], s[231:224], s[223:216], s[215:208], s[207:200], s[199:192]};
	a[0][4] = {s[319:312], s[311:304], s[303:296], s[295:288], s[287:280], s[279:272], s[271:264], s[263:256]};
	
	a[1][0] = {s[383:376], s[375:368], s[367:360], s[359:352], s[351:344], s[343:336], s[335:328], s[327:320]};
	a[1][1] = {s[447:440], s[439:432], s[431:424], s[423:416], s[415:408], s[407:400], s[399:392], s[391:384]};
	a[1][2] = {s[511:504], s[503:496], s[495:488], s[487:480], s[479:472], s[471:464], s[463:456], s[455:448]};
	a[1][3] = {s[575:568], s[567:560], s[559:552], s[551:544], s[543:536], s[535:528], s[527:520], s[519:512]};
	a[1][4] = {s[639:632], s[631:624], s[623:616], s[615:608], s[607:600], s[599:592], s[591:584], s[583:576]};

	a[2][0] = {s[703:696], s[695:688], s[687:680], s[679:672], s[671:664], s[663:656], s[655:648], s[647:640]};
	a[2][1] = {s[767:760], s[759:752], s[751:744], s[743:736], s[735:728], s[727:720], s[719:712], s[711:704]};
	a[2][2] = {s[831:824], s[823:816], s[815:808], s[807:800], s[799:792], s[791:784], s[783:776], s[775:768]};
	a[2][3] = {s[895:888], s[887:880], s[879:872], s[871:864], s[863:856], s[855:848], s[847:840], s[839:832]};
	a[2][4] = {s[959:952], s[951:944], s[943:936], s[935:928], s[927:920], s[919:912], s[911:904], s[903:896]};

	a[3][0] = {s[1023:1016], s[1015:1008], s[1007:1000], s[999:992], s[991:984], s[983:976], s[975:968], s[967:960]};
	a[3][1] = {s[1087:1080], s[1079:1072], s[1071:1064], s[1063:1056], s[1055:1048], s[1047:1040], s[1039:1032], s[1031:1024]};
	a[3][2] = {s[1151:1144], s[1143:1136], s[1135:1128], s[1127:1120], s[1119:1112], s[1111:1104], s[1103:1096], s[1095:1088]};
	a[3][3] = {s[1215:1208], s[1207:1200], s[1199:1192], s[1191:1184], s[1183:1176], s[1175:1168], s[1167:1160], s[1159:1152]};
	a[3][4] = {s[1279:1272], s[1271:1264], s[1264:1256], s[1255:1248], s[1247:1240], s[1239:1232], s[1231:1224], s[1223:1216]};

	a[4][0] = {s[1343:1336], s[1335:1328], s[1327:1320], s[1319:1312], s[1311:1304], s[1303:1296], s[1295:1288], s[1287:1280]};
	a[4][1] = {s[1407:1400], s[1399:1392], s[1391:1384], s[1383:1376], s[1375:1368], s[1367:1360], s[1359:1352], s[1351:1344]};
	a[4][2] = {s[1471:1464], s[1463:1456], s[1455:1448], s[1447:1440], s[1439:1432], s[1431:1424], s[1423:1416], s[1415:1408]};
	a[4][3] = {s[1535:1528], s[1527:1520], s[1519:1512], s[1511:1504], s[1503:1496], s[1495:1488], s[1487:1480], s[1479:1472]};
	a[4][4] = {s[1599:1592], s[1591:1584], s[1583:1576], s[1575:1568], s[1567:1560], s[1559:1552], s[1551:1544], s[1543:1536]};
	*/
	a[0][0] = s[63:0];
	a[0][1] = s[127:64]; 
	a[0][2] = s[191:128];
	a[0][3] = s[255:192];
	a[0][4] = s[319:256];

	a[1][0] = s[383:320];
	a[1][1] = s[447:384];
	a[1][2] = s[511:448];
	a[1][3] = s[575:512];
	a[1][4] = s[639:576];
	
	a[2][0] = s[703:640];
	a[2][1] = s[767:704];
	a[2][2] = s[831:768];
	a[2][3] = s[895:832];
	a[2][4] = s[959:896];

	a[3][0] = s[1023:960];
	a[3][1] = s[1087:1024];
	a[3][2] = s[1151:1088];
	a[3][3] = s[1215:1152];
	a[3][4] = s[1279:1216];
	
	a[4][0] = s[1343:1280];
	a[4][1] = s[1407:1344];
	a[4][2] = s[1471:1408];
	a[4][3] = s[1535:1472];
	a[4][4] = s[1599:1536];
	
end	
endmodule

module string_to_array_tb();
logic		[1599:0] init_state;
logic   	[1343:0] data_in;
logic 		[2:0]	 c_mode;
logic		[1599:0] s;
state a;

VSX_module VSX(data_in, init_state, c_mode, s);
string_to_array sta(s,a);

initial 
begin
//s = 1600'h0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef_0123_4567_89ab_cdef;
data_in = 1344'h000000000000000000000000000000000000000000000000000000000000000080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000600000000000000000000000000000000;
init_state = 0;
c_mode = 1;
#5;
end

endmodule